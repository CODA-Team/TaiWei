# BSD 3-Clause License
# 
# Copyright 2020 Lawrence T. Clark, Vinay Vashishtha, or Arizona State
# University
# 
# Redistribution and use in source and binary forms, with or without
# modification, are permitted provided that the following conditions are met:
# 
# 1. Redistributions of source code must retain the above copyright notice,
# this list of conditions and the following disclaimer.
# 
# 2. Redistributions in binary form must reproduce the above copyright
# notice, this list of conditions and the following disclaimer in the
# documentation and/or other materials provided with the distribution.
# 
# 3. Neither the name of the copyright holder nor the names of its
# contributors may be used to endorse or promote products derived from this
# software without specific prior written permission.
# 
# THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
# AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
# IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
# ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
# LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
# CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
# SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
# INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
# CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
# ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
# POSSIBILITY OF SUCH DAMAGE.

VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
CLEARANCEMEASURE EUCLIDEAN ;
USEMINSPACING OBS OFF ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.001 ;

# ========================
# Property Definitions
# ========================
PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_PITCH STRING ;
  LAYER LEF58_GAP STRING ;
  LAYER LEF58_EOLKEEPOUT STRING ;
  LAYER LEF58_SPACING STRING ;
  LAYER LEF58_CORNERSPACING STRING ;
  LAYER LEF58_WIDTHTABLE STRING ;
  LAYER LEF58_CUTCLASS STRING ;
  LAYER LEF58_SPACINGTABLE STRING ;
  LAYER LEF58_ENCLOSURE STRING ;
  LAYER LEF58_RIGHTWAYONGRIDONLY STRING ;
  LAYER LEF58_RECTONLY STRING ;
END PROPERTYDEFINITIONS

# ======================================================
# 1) LAYER DEFINITIONS (all layers first, ordered)
# ======================================================

# --- Base / Implants / Wells ---
LAYER LVTN
  TYPE IMPLANT ;
END LVTN

LAYER LVTP
  TYPE IMPLANT ;
END LVTP

LAYER RVTN
  TYPE IMPLANT ;
END RVTN

LAYER RVTP
  TYPE IMPLANT ;
END RVTP

LAYER RVTN_m
  TYPE IMPLANT ;
END RVTN_m

LAYER RVTP_m
  TYPE IMPLANT ;
END RVTP_m

LAYER SLVTN
  TYPE IMPLANT ;
END SLVTN

LAYER SLVTP
  TYPE IMPLANT ;
END SLVTP

LAYER nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END pwell

LAYER Gate
  TYPE MASTERSLICE ;
END Gate

LAYER Active
  TYPE MASTERSLICE ;
END Active

# --- Bottom die stack (bottom-up) ---
# LAYER V0
#   TYPE CUT ;
#   SPACING 0.018 ;
#   WIDTH 0.018 ;
# END V0

LAYER M1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.036 ;
  WIDTH 0.018 ;
  SPACING 0.018 ;
  AREA 0.000666 ;
  SPACING 0.018 RANGE 0.036 1.0 ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.01825 EXTENSION 0.0 0.0 0.031 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERONLY 0.01 WIDTH 0.018 SPACING 0.018 ;" ;
  OFFSET 0.0 ;
# --- RC added from ict/setRC for M1 ---
  THICKNESS 0.036 ;
  HEIGHT 0.141 ;
  RESISTANCE RPERSQ 1.267515 ;
  CAPACITANCE CPERSQDIST 1.000000e-08 ;
  EDGECAPACITANCE 1.000000e-08 ;
END M1

LAYER V1
  TYPE CUT ;
  SPACING 0.018 ;
  WIDTH 0.018 ;
# --- RC added from ict/setRC for V1 ---
  RESISTANCE 17.2 ;
END V1

LAYER M2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.018 ;
  SPACING 0.018 ;
  OFFSET -0.27 ;
  AREA 0.000666 ;
  MINSIZE 0.037 0.018 ;
  PITCH 0.045 0.036 ;
  PROPERTY LEF58_PITCH "
   PITCH 0.036 FIRSTLASTPITCH 0.045
     ;
   " ;
  PROPERTY LEF58_SPACING
   " SPACING 0.018 ENDOFLINE 0.025 WITHIN 0.02 ENDTOEND 0.031
     PARALLELEDGE 0.025 WITHIN 0.02 ; " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.025 EXTENSION 0.0 0.0125 0.031 CORNERONLY ;
   " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER WIDTH 0.0 SPACING 0.02 ;
   " ;
  PROPERTY LEF58_WIDTHTABLE "
   WIDTHTABLE 0.018 0.09 0.162 0.234 0.306 0.378 ;
   " ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M2 ---
  THICKNESS 0.036 ;
  HEIGHT 0.213 ;
  RESISTANCE RPERSQ 0.83216 ;
  CAPACITANCE CPERSQDIST 0.003076 ;
  EDGECAPACITANCE 6.458970e-05 ;
END M2

LAYER V2
  TYPE CUT ;
  SPACING 0.018 ;
  WIDTH 0.018 ;
# --- RC added from ict/setRC for V2 ---
  RESISTANCE 17.2 ;
END V2

LAYER M3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.036 ;
  OFFSET 0.0 ;
  WIDTH 0.018 ;
  SPACING 0.018 ;
  AREA 0.000666 ;
  MINSIZE 0.037 0.018 ;
  PROPERTY LEF58_SPACING
   " SPACING 0.018 ENDOFLINE 0.025 WITHIN 0.0125 ENDTOEND 0.031
     PARALLELEDGE 0.025 WITHIN 0.02 ; " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.025 EXTENSION 0.0 0.0125 0.031 CORNERONLY ;
   " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER WIDTH 0.0 SPACING 0.02 ;
   " ;
  PROPERTY LEF58_WIDTHTABLE
   " WIDTHTABLE 0.018 0.09 0.162 0.234 0.306 0.378 ; " ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M3 ---
  THICKNESS 0.036 ;
  HEIGHT 0.285 ;
  RESISTANCE RPERSQ 0.653852 ;
  CAPACITANCE CPERSQDIST 0.002566 ;
  EDGECAPACITANCE 5.388425e-05 ;
END M3

LAYER V3
  TYPE CUT ;
  PROPERTY LEF58_CUTCLASS "
   CUTCLASS V3 WIDTH 0.018 LENGTH 0.024 CUTS 1 ;
   CUTCLASS V3_0p480 WIDTH 0.018 LENGTH 0.12 CUTS 4 ;
   CUTCLASS V3_0p864 WIDTH 0.018 LENGTH 0.216 CUTS 8 ;
   " ;
  PROPERTY LEF58_SPACINGTABLE "
      SPACINGTABLE
       DEFAULT 0.034
       CUTCLASS V3 V3_0p480 V3_0p864
              V3       -  -        -        -  - -
              V3_0p480 -  -        -        -  - -
              V3_0p864 -  -        -        -  - -
      ;
   " ;
  PROPERTY LEF58_ENCLOSURE "
   ENCLOSURE CUTCLASS V3 BELOW EOL 0.0 0.005 0.0 ;
   ENCLOSURE CUTCLASS V3 ABOVE EOL 0.02425 0.011 0.0 ;
   ENCLOSURE CUTCLASS V3_0p480 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS V3_0p864 END 0.0 SIDE 0.0 ;
   " ;
# --- RC added from ict/setRC for V3 ---
  RESISTANCE 17.2 ;
END V3

LAYER M4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.048 ;
  WIDTH 0.024 ;
  SPACING 0.024 ;
  OFFSET 0.003 ;
  AREA 0.002 ;
  PROPERTY LEF58_SPACING " SPACING 0.024 ENDOFLINE 0.025 WITHIN 0.04 ENDTOEND 0.04 ; " ;
  PROPERTY LEF58_WIDTHTABLE " WIDTHTABLE 0.024 0.12 0.216 0.312 0.408 ; " ;
  PROPERTY LEF58_CORNERSPACING "   CORNERSPACING CONVEXCORNER CORNERONLY 0.048
   WIDTH 0.0 SPACING 0.04 ;
   " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.025 EXTENSION 0.048 0.02425 0.048 CORNERONLY ;
   " ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0
    WIDTH 0.0 0.024
    WIDTH 0.025 0.072 ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M4 ---
  THICKNESS 0.048 ;
  HEIGHT 0.357 ;
  RESISTANCE RPERSQ 0.487399 ;
  CAPACITANCE CPERSQDIST 0.002368 ;
  EDGECAPACITANCE 6.630190e-05 ;
END M4

LAYER V4
  TYPE CUT ;
  PROPERTY LEF58_CUTCLASS "
   CUTCLASS Vx WIDTH 0.024 LENGTH 0.024 ;
   CUTCLASS Vx_0p480 WIDTH 0.024 LENGTH 0.12 CUTS 4 ;
   CUTCLASS Vx_0p864 WIDTH 0.024 LENGTH 0.216 CUTS 8 ;
   CUTCLASS Vx_1p248 WIDTH 0.024 LENGTH 0.312 CUTS 12 ;
   CUTCLASS Vx_1p632 WIDTH 0.024 LENGTH 0.408 CUTS 16 ;
   " ;
  PROPERTY LEF58_SPACINGTABLE "
      SPACINGTABLE
       DEFAULT 0.034
       CUTCLASS Vx Vx_0p480 Vx_0p864 Vx_1p248 Vx_1p632
              Vx       -  -        -        -        - -  -        -        -        -
              Vx_0p480 -  -        -        -        - -  -        -        -        -
	      Vx_0p864 -  -        -        -        - -  -        -        -        -
	      Vx_1p248 -  -        -        -        - -  -        -        -        -
	      Vx_1p632 -  -        -        -        - -  -        -        -        -
      ;
   " ;
  PROPERTY LEF58_ENCLOSURE "
   ENCLOSURE CUTCLASS Vx 0.011 0.0 ;
   ENCLOSURE CUTCLASS Vx EOL 0.0 0.011 0.011 ;
   ENCLOSURE CUTCLASS Vx_0p480 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_0p864 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p248 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p632 END 0.0 SIDE 0.0 ;
   " ;
# --- RC added from ict/setRC for V4 ---
  RESISTANCE 11.8 ;
END V4

LAYER M5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.048 ;
  WIDTH 0.024 ;
  SPACING 0.024 ;
  OFFSET 0.0 ;
  AREA 0.002 ;
  PROPERTY LEF58_SPACING " SPACING 0.024 ENDOFLINE 0.025 WITHIN 0.04 ENDTOEND 0.04 ; " ;
  MINIMUMDENSITY 15.0 ;
  MAXIMUMDENSITY 90.0 ;
  DENSITYCHECKWINDOW 20.0 20.0 ;
  DENSITYCHECKSTEP 10.0 ;
  PROPERTY LEF58_WIDTHTABLE
   " WIDTHTABLE 0.024 0.12 0.216 0.312 0.408 0.504 0.6 0.696 0.792 0.888 0.984 ; " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER CORNERONLY 0.048
   WIDTH 0.0 SPACING 0.04 ;
   " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.025 EXTENSION 0.048 0.02425 0.048
      CORNERONLY ;
   " ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0
    WIDTH 0.0 0.024
    WIDTH 0.025 0.072 ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M5 ---
  THICKNESS 0.048 ;
  HEIGHT 0.453 ;
  RESISTANCE RPERSQ 0.463212 ;
  CAPACITANCE CPERSQDIST 0.002145 ;
  EDGECAPACITANCE 6.005755e-05 ;
END M5

LAYER V5
  TYPE CUT ;
  PROPERTY LEF58_CUTCLASS "
   CUTCLASS Vx WIDTH 0.024 LENGTH 0.032 ;
   CUTCLASS Vx_0p480 WIDTH 0.024 LENGTH 0.16 CUTS 4 ;
   CUTCLASS Vx_0p864 WIDTH 0.024 LENGTH 0.288 CUTS 8 ;
   CUTCLASS Vx_1p248 WIDTH 0.024 LENGTH 0.416 CUTS 12 ;
   CUTCLASS Vx_1p632 WIDTH 0.024 LENGTH 0.544 CUTS 16 ;
   " ;
  PROPERTY LEF58_SPACINGTABLE "
      SPACINGTABLE
       DEFAULT 0.034
       CUTCLASS Vx Vx_0p480 Vx_0p864 Vx_1p248 Vx_1p632
              Vx       -  -        -        -        - -  -        -        -        -
              Vx_0p480 -  -        -        -        - -  -        -        -        -
	      Vx_0p864 -  -        -        -        - -  -        -        -        -
	      Vx_1p248 -  -        -        -        - -  -        -        -        -
	      Vx_1p632 -  -        -        -        - -  -        -        -        -
      ;
   " ;
  PROPERTY LEF58_ENCLOSURE "
   ENCLOSURE CUTCLASS Vx EOL 0.02425 0.011 0.011 ;
   ENCLOSURE CUTCLASS Vx_0p480 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_0p864 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p248 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p632 END 0.0 SIDE 0.0 ;
   " ;
# --- RC added from ict/setRC for V5 ---
  RESISTANCE 11.8 ;
END V5

LAYER M6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.064 ;
  WIDTH 0.032 ;
  SPACING 0.032 ;
  AREA 0.0021875 ;
  PROPERTY LEF58_SPACING
   " SPACING 0.032 ENDOFLINE 0.0375 WITHIN 0.04 ENDTOEND 0.04 ; " ;
  PROPERTY LEF58_WIDTHTABLE " WIDTHTABLE 0.032 0.16 0.288 0.416 0.544 ; " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER CORNERONLY 0.048
   WIDTH 0.0 SPACING 0.04 ;
   " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.05 EXTENSION 0.048 0.03225 0.048 CORNERONLY ;
   " ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0
    WIDTH 0.0 0.032
    WIDTH 0.033 0.072 ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M6 ---
  THICKNESS 0.064 ;
  HEIGHT 0.549 ;
  RESISTANCE RPERSQ 0.379581 ;
  CAPACITANCE CPERSQDIST 0.001651 ;
  EDGECAPACITANCE 6.165110e-05 ;
END M6

LAYER V6
  TYPE CUT ;
  PROPERTY LEF58_CUTCLASS "
   CUTCLASS Vx WIDTH 0.032 LENGTH 0.032 ;
   CUTCLASS Vx_0p640 WIDTH 0.032 LENGTH 0.16 CUTS 4 ;
   CUTCLASS Vx_1p152 WIDTH 0.032 LENGTH 0.288 CUTS 8 ;
   CUTCLASS Vx_1p664 WIDTH 0.032 LENGTH 0.416 CUTS 12 ;
   CUTCLASS Vx_2p176 WIDTH 0.032 LENGTH 0.544 CUTS 16 ;
   " ;
  PROPERTY LEF58_SPACINGTABLE "
      SPACINGTABLE
       DEFAULT 0.034
       CUTCLASS Vx Vx_0p640 Vx_1p152 Vx_1p664 Vx_2p176
              Vx       -  -        -        -        - -  -        -        -        -
              Vx_0p640 -  -        -        -        - -  -        -        -        -
	      Vx_1p152 -  -        -        -        - -  -        -        -        -
	      Vx_1p664 -  -        -        -        - -  -        -        -        -
	      Vx_2p176 -  -        -        -        - -  -        -        -        -
      ;
   " ;
  PROPERTY LEF58_ENCLOSURE "
   ENCLOSURE CUTCLASS Vx 0.011 0.0 ;
   ENCLOSURE CUTCLASS Vx EOL 0.0 0.011 0.011 ;
   ENCLOSURE CUTCLASS Vx_0p640 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p152 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p664 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_2p176 END 0.0 SIDE 0.0 ;
   " ;
# --- RC added from ict/setRC for V6 ---
  RESISTANCE 8.2 ;
END V6

LAYER M7
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.064 ;
  WIDTH 0.032 ;
  SPACING 0.032 ;
  AREA 0.0021875 ;
  PROPERTY LEF58_SPACING
   " SPACING 0.03 ENDOFLINE 0.0375 WITHIN 0.04 ENDTOEND 0.04 ; " ;
  PROPERTY LEF58_WIDTHTABLE " WIDTHTABLE 0.032 0.16 0.288 0.416 0.544 ; " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER CORNERONLY 0.075
   WIDTH 0.0 SPACING 0.04 ;
   " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.05 EXTENSION 0.048 0.03225 0.048
      CORNERONLY ;
   " ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0
    WIDTH 0.0 0.032
    WIDTH 0.033 0.072 ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M7 ---
  THICKNESS 0.064 ;
  HEIGHT 0.677 ;
  RESISTANCE RPERSQ 0.400995 ;
  CAPACITANCE CPERSQDIST 0.001378 ;
  EDGECAPACITANCE 5.146050e-05 ;
END M7

LAYER hb_layer
  TYPE CUT ;
  SPACING 0.5 ;
  WIDTH 0.5 ;
  RESISTANCE 0.02 ;
END hb_layer

LAYER M6_m
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.064 ;
  WIDTH 0.032 ;
  SPACING 0.032 ;
  AREA 0.0021875 ;
  PROPERTY LEF58_SPACING " SPACING 0.032 ENDOFLINE 0.0375 WITHIN 0.04 ENDTOEND 0.04 ; " ;
  PROPERTY LEF58_WIDTHTABLE " WIDTHTABLE 0.032 0.16 0.288 0.416 0.544 ; " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER CORNERONLY 0.048
   WIDTH 0.0 SPACING 0.04 ;
   " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.05 EXTENSION 0.048 0.03225 0.048 CORNERONLY ;
   " ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0
    WIDTH 0.0 0.032
    WIDTH 0.033 0.072 ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M6_m ---
  THICKNESS 0.064 ;
  HEIGHT 1.701 ;
  RESISTANCE RPERSQ 0.379581 ;
  CAPACITANCE CPERSQDIST 0.001651 ;
  EDGECAPACITANCE 6.165110e-05 ;
END M6_m

LAYER V5_m
  TYPE CUT ;
  PROPERTY LEF58_CUTCLASS "
   CUTCLASS Vx WIDTH 0.024 LENGTH 0.032 ;
   CUTCLASS Vx_0p480 WIDTH 0.024 LENGTH 0.16 CUTS 4 ;
   CUTCLASS Vx_0p864 WIDTH 0.024 LENGTH 0.288 CUTS 8 ;
   CUTCLASS Vx_1p248 WIDTH 0.024 LENGTH 0.416 CUTS 12 ;
   CUTCLASS Vx_1p632 WIDTH 0.024 LENGTH 0.544 CUTS 16 ;
   " ;
  PROPERTY LEF58_SPACINGTABLE "
      SPACINGTABLE
       DEFAULT 0.034
       CUTCLASS Vx Vx_0p480 Vx_0p864 Vx_1p248 Vx_1p632
              Vx       -  -        -        -        - -  -        -        -        -
              Vx_0p480 -  -        -        -        - -  -        -        -        -
	      Vx_0p864 -  -        -        -        - -  -        -        -        -
	      Vx_1p248 -  -        -        -        - -  -        -        -        -
	      Vx_1p632 -  -        -        -        - -  -        -        -        -
      ;
   " ;
  PROPERTY LEF58_ENCLOSURE "
   ENCLOSURE CUTCLASS Vx EOL 0.02425 0.011 0.011 ;
   ENCLOSURE CUTCLASS Vx_0p480 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_0p864 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p248 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p632 END 0.0 SIDE 0.0 ;
   " ;
# --- RC added from ict/setRC for V5_m ---
  RESISTANCE 11.8 ;
END V5_m

LAYER M5_m
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.048 ;
  WIDTH 0.024 ;
  SPACING 0.024 ;
  OFFSET 0.0 ;
  AREA 0.002 ;
  PROPERTY LEF58_SPACING " SPACING 0.024 ENDOFLINE 0.025 WITHIN 0.04 ENDTOEND 0.04 ; " ;
  MINIMUMDENSITY 15.0 ;
  MAXIMUMDENSITY 90.0 ;
  DENSITYCHECKWINDOW 20.0 20.0 ;
  DENSITYCHECKSTEP 10.0 ;
  PROPERTY LEF58_WIDTHTABLE
   " WIDTHTABLE 0.024 0.12 0.216 0.312 0.408 0.504 0.6 0.696 0.792 0.888 0.984 ; " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER CORNERONLY 0.048
   WIDTH 0.0 SPACING 0.04 ;
   " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.025 EXTENSION 0.048 0.02425 0.048
      CORNERONLY ;
   " ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0
    WIDTH 0.0 0.024
    WIDTH 0.025 0.072 ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M5_m ---
  THICKNESS 0.048 ;
  HEIGHT 1.797 ;
  RESISTANCE RPERSQ 0.463212 ;
  CAPACITANCE CPERSQDIST 0.002145 ;
  EDGECAPACITANCE 6.005755e-05 ;
END M5_m

LAYER V4_m
  TYPE CUT ;
  PROPERTY LEF58_CUTCLASS "
   CUTCLASS Vx WIDTH 0.024 LENGTH 0.024 ;
   CUTCLASS Vx_0p480 WIDTH 0.024 LENGTH 0.12 CUTS 4 ;
   CUTCLASS Vx_0p864 WIDTH 0.024 LENGTH 0.216 CUTS 8 ;
   CUTCLASS Vx_1p248 WIDTH 0.024 LENGTH 0.312 CUTS 12 ;
   CUTCLASS Vx_1p632 WIDTH 0.024 LENGTH 0.408 CUTS 16 ;
   " ;
  PROPERTY LEF58_SPACINGTABLE "
      SPACINGTABLE
       DEFAULT 0.034
       CUTCLASS Vx Vx_0p480 Vx_0p864 Vx_1p248 Vx_1p632
              Vx       -  -        -        -        - -  -        -        -        -
              Vx_0p480 -  -        -        -        - -  -        -        -        -
	      Vx_0p864 -  -        -        -        - -  -        -        -        -
	      Vx_1p248 -  -        -        -        - -  -        -        -        -
	      Vx_1p632 -  -        -        -        - -  -        -        -        -
      ;
   " ;
  PROPERTY LEF58_ENCLOSURE "
   ENCLOSURE CUTCLASS Vx 0.011 0.0 ;
   ENCLOSURE CUTCLASS Vx EOL 0.0 0.011 0.011 ;
   ENCLOSURE CUTCLASS Vx_0p480 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_0p864 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p248 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p632 END 0.0 SIDE 0.0 ;
   " ;
# --- RC added from ict/setRC for V4_m ---
  RESISTANCE 11.8 ;
END V4_m

LAYER M4_m
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.048 ;
  WIDTH 0.024 ;
  SPACING 0.024 ;
  OFFSET 0.003 ;
  AREA 0.002 ;
  PROPERTY LEF58_SPACING " SPACING 0.024 ENDOFLINE 0.025 WITHIN 0.04 ENDTOEND 0.04 ; " ;
  PROPERTY LEF58_WIDTHTABLE " WIDTHTABLE 0.024 0.12 0.216 0.312 0.408 ; " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER CORNERONLY 0.048
   WIDTH 0.0 SPACING 0.04 ;
   " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.025 EXTENSION 0.048 0.02425 0.048 CORNERONLY ;
   " ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0
    WIDTH 0.0 0.024
    WIDTH 0.025 0.072 ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M4_m ---
  THICKNESS 0.048 ;
  HEIGHT 1.893 ;
  RESISTANCE RPERSQ 0.487399 ;
  CAPACITANCE CPERSQDIST 0.002368 ;
  EDGECAPACITANCE 6.630190e-05 ;
END M4_m

LAYER V3_m
  TYPE CUT ;
  PROPERTY LEF58_CUTCLASS "
   CUTCLASS V3 WIDTH 0.018 LENGTH 0.024 CUTS 1 ;
   CUTCLASS V3_0p480 WIDTH 0.018 LENGTH 0.12 CUTS 4 ;
   CUTCLASS V3_0p864 WIDTH 0.018 LENGTH 0.216 CUTS 8 ;
   " ;
  PROPERTY LEF58_SPACINGTABLE "
      SPACINGTABLE
       DEFAULT 0.034
       CUTCLASS V3 V3_0p480 V3_0p864
              V3       -  -        -        -  - -
              V3_0p480 -  -        -        -  - -
              V3_0p864 -  -        -        -  - -
      ;
   " ;
  PROPERTY LEF58_ENCLOSURE "
   ENCLOSURE CUTCLASS V3 BELOW EOL 0.0 0.005 0.0 ;
   ENCLOSURE CUTCLASS V3 ABOVE EOL 0.02425 0.011 0.0 ;
   ENCLOSURE CUTCLASS V3_0p480 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS V3_0p864 END 0.0 SIDE 0.0 ;
   " ;
# --- RC added from ict/setRC for V3_m ---
  RESISTANCE 17.2 ;
END V3_m

LAYER M3_m
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.036 ;
  OFFSET 0.0 ;
  WIDTH 0.018 ;
  SPACING 0.018 ;
  AREA 0.000666 ;
  MINSIZE 0.037 0.018 ;
  PROPERTY LEF58_SPACING
   " SPACING 0.018 ENDOFLINE 0.025 WITHIN 0.0125 ENDTOEND 0.031
     PARALLELEDGE 0.025 WITHIN 0.02 ; " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.025 EXTENSION 0.0 0.0125 0.031 CORNERONLY ;
   " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER WIDTH 0.0 SPACING 0.02
     ;
   " ;
  PROPERTY LEF58_WIDTHTABLE
   " WIDTHTABLE 0.018 0.09 0.162 0.234 0.306 0.378 ; " ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M3_m ---
  THICKNESS 0.036 ;
  HEIGHT 1.965 ;
  RESISTANCE RPERSQ 0.653852 ;
  CAPACITANCE CPERSQDIST 0.002566 ;
  EDGECAPACITANCE 5.388425e-05 ;
END M3_m

LAYER V2_m
  TYPE CUT ;
  SPACING 0.018 ;
  WIDTH 0.018 ;
# --- RC added from ict/setRC for V2_m ---
  RESISTANCE 17.2 ;
END V2_m

LAYER M2_m
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.018 ;
  SPACING 0.018 ;
  OFFSET -0.27 ;
  AREA 0.000666 ;
  MINSIZE 0.037 0.018 ;
  PITCH 0.045 0.036 ;
  PROPERTY LEF58_PITCH "
   PITCH 0.036 FIRSTLASTPITCH 0.045
     ;
   " ;
  PROPERTY LEF58_SPACING
   " SPACING 0.018 ENDOFLINE 0.025 WITHIN 0.02 ENDTOEND 0.031
     PARALLELEDGE 0.025 WITHIN 0.02 ; " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.025 EXTENSION 0.0 0.0125 0.031 CORNERONLY ;
   " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER WIDTH 0.0 SPACING 0.02 ;
   " ;
  PROPERTY LEF58_WIDTHTABLE "
   WIDTHTABLE 0.018 0.09 0.162 0.234 0.306 0.378 ;
   " ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M2_m ---
  THICKNESS 0.036 ;
  HEIGHT 2.037 ;
  RESISTANCE RPERSQ 0.83216 ;
  CAPACITANCE CPERSQDIST 0.003076 ;
  EDGECAPACITANCE 6.458970e-05 ;
END M2_m

LAYER V1_m
  TYPE CUT ;
  SPACING 0.018 ;
  WIDTH 0.018 ;
# --- RC added from ict/setRC for V1_m ---
  RESISTANCE 17.2 ;
END V1_m

LAYER M1_m
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.036 ;
  WIDTH 0.018 ;
  SPACING 0.018 ;
  AREA 0.000666 ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.01825 EXTENSION 0.0 0.0 0.031 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERONLY 0.01 WIDTH 0.018 SPACING 0.018 ;" ;
  OFFSET 0.0 ;
# --- RC added from ict/setRC for M1_m ---
  THICKNESS 0.036 ;
  HEIGHT 2.109 ;
  RESISTANCE RPERSQ 1.267515 ;
  CAPACITANCE CPERSQDIST 1.000000e-08 ;
  EDGECAPACITANCE 1.000000e-08 ;
END M1_m

# LAYER V0_m
#   TYPE CUT ;
#   SPACING 0.018 ;
#   WIDTH 0.018 ;
# END V0_m
LAYER V1_add
  TYPE CUT ;
  SPACING 0.018 ;
  WIDTH 0.018 ;
# --- RC added from ict/setRC for V1_add ---
  RESISTANCE 17.2 ;
END V1_add

LAYER M2_add
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.018 ;
  SPACING 0.018 ;
  OFFSET -0.27 ;
  AREA 0.000666 ;
  MINSIZE 0.037 0.018 ;
  PITCH 0.045 0.036 ;
  PROPERTY LEF58_PITCH "
   PITCH 0.036 FIRSTLASTPITCH 0.045
     ;
  " ;
  PROPERTY LEF58_SPACING
   " SPACING 0.018 ENDOFLINE 0.025 WITHIN 0.02 ENDTOEND 0.031
     PARALLELEDGE 0.025 WITHIN 0.02 ; " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.025 EXTENSION 0.0 0.0125 0.031 CORNERONLY ;
  " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER WIDTH 0.0 SPACING 0.02 ;
  " ;
  PROPERTY LEF58_WIDTHTABLE "
   WIDTHTABLE 0.018 0.09 0.162 0.234 0.306 0.378 ;
  " ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY "
    RIGHTWAYONGRIDONLY ;
  " ;
  PROPERTY LEF58_RECTONLY "
    RECTONLY ;
  " ;
# --- RC added from ict/setRC for M2_add ---
  THICKNESS 0.036 ;
  HEIGHT 2.181 ;
  RESISTANCE RPERSQ 0.83216 ;
  CAPACITANCE CPERSQDIST 0.003076 ;
  EDGECAPACITANCE 6.458970e-05 ;
END M2_add

LAYER V2_add
  TYPE CUT ;
  SPACING 0.018 ;
  WIDTH 0.018 ;
# --- RC added from ict/setRC for V2_add ---
  RESISTANCE 17.2 ;
END V2_add

LAYER M3_add
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.036 ;
  OFFSET 0.0 ;
  WIDTH 0.018 ;
  SPACING 0.018 ;
  AREA 0.000666 ;
  MINSIZE 0.037 0.018 ;
  PROPERTY LEF58_SPACING
   " SPACING 0.018 ENDOFLINE 0.025 WITHIN 0.0125 ENDTOEND 0.031
     PARALLELEDGE 0.025 WITHIN 0.02 ; " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.025 EXTENSION 0.0 0.0125 0.031 CORNERONLY ;
  " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER WIDTH 0.0 SPACING 0.02 ;
  " ;
  PROPERTY LEF58_WIDTHTABLE
   " WIDTHTABLE 0.018 0.09 0.162 0.234 0.306 0.378 ; " ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY "
    RIGHTWAYONGRIDONLY ;
  " ;
  PROPERTY LEF58_RECTONLY "
    RECTONLY ;
  " ;
# --- RC added from ict/setRC for M3_add ---
  THICKNESS 0.036 ;
  HEIGHT 2.253 ;
  RESISTANCE RPERSQ 0.653852 ;
  CAPACITANCE CPERSQDIST 0.002566 ;
  EDGECAPACITANCE 5.388425e-05 ;
END M3_add

VIA VIA12 Default
  LAYER M1 ;  RECT -0.009 -0.011 0.009 0.011 ;
  LAYER M2 ;  RECT -0.014 -0.009 0.014 0.009 ;
  LAYER V1 ;  RECT -0.009 -0.009 0.009 0.009 ;
END VIA12

VIA VIA23 Default
  LAYER M2 ;  RECT -0.014 -0.009 0.014 0.009 ;
  LAYER M3 ;  RECT -0.009 -0.014 0.009 0.014 ;
  LAYER V2 ;  RECT -0.009 -0.009 0.009 0.009 ;
END VIA23

VIA VIA34 Default
  LAYER M3 ;  RECT -0.009 -0.017 0.009 0.017 ;
  LAYER M4 ;  RECT -0.02 -0.012 0.02 0.012 ;
  LAYER V3 ;  RECT -0.009 -0.012 0.009 0.012 ;
END VIA34

VIA VIA45 Default
  LAYER M4 ;  RECT -0.023 -0.012 0.023 0.012 ;
  LAYER M5 ;  RECT -0.012 -0.023 0.012 0.023 ;
  LAYER V4 ;  RECT -0.012 -0.012 0.012 0.012 ;
END VIA45

VIA VIA56 Default
  LAYER M5 ;  RECT -0.012 -0.027 0.012 0.027 ;
  LAYER M6 ;  RECT -0.023 -0.016 0.023 0.016 ;
  LAYER V5 ;  RECT -0.012 -0.016 0.012 0.016 ;
END VIA56

VIA VIA67 Default
  LAYER M6 ;  RECT -0.027 -0.016 0.027 0.016 ;
  LAYER M7 ;  RECT -0.016 -0.027 0.016 0.027 ;
  LAYER V6 ;  RECT -0.016 -0.016 0.016 0.016 ;
END VIA67

VIA hb_layer_0 DEFAULT
  LAYER hb_layer ; RECT -0.25 -0.25 0.25 0.25 ;
  LAYER M7 ; RECT -0.25 -0.25 0.25 0.25 ;
  LAYER M6_m ; RECT -0.25 -0.25 0.25 0.25 ;
END hb_layer_0
VIA hb_layer_1 DEFAULT
  LAYER hb_layer ; RECT -0.25 -0.25 0.25 0.25 ;
  LAYER M7 ; RECT -0.5 -0.5 0.5 0.5 ;
  LAYER M6_m ; RECT -0.25 -0.5 0.25 0.5 ;
END hb_layer_1
VIA hb_layer_2 DEFAULT
  LAYER hb_layer ; RECT -0.25 -0.25 0.25 0.25 ;
  LAYER M7 ; RECT -0.5 -0.5 0.5 0.5 ;
  LAYER M6_m ; RECT -0.5 -0.25 0.5 0.25 ;
END hb_layer_2
VIA hb_layer_3 DEFAULT
  LAYER hb_layer ; RECT -0.25 -0.25 0.25 0.25 ;
  LAYER M7 ; RECT -0.25 -0.5 0.25 0.5 ;
  LAYER M6_m ; RECT -0.5 -0.5 0.5 0.5 ;
END hb_layer_3
VIA hb_layer_4 DEFAULT
  LAYER hb_layer ; RECT -0.25 -0.25 0.25 0.25 ;
  LAYER M7 ; RECT -0.25 -0.5 0.25 0.5 ;
  LAYER M6_m ; RECT -0.25 -0.5 0.25 0.5 ;
END hb_layer_4
VIA hb_layer_5 DEFAULT
  LAYER hb_layer ; RECT -0.25 -0.25 0.25 0.25 ;
  LAYER M7 ; RECT -0.25 -0.5 0.25 0.5 ;
  LAYER M6_m ; RECT -0.5 -0.25 0.5 0.25 ;
END hb_layer_5
VIA hb_layer_6 DEFAULT
  LAYER hb_layer ; RECT -0.25 -0.25 0.25 0.25 ;
  LAYER M7 ; RECT -0.5 -0.25 0.5 0.25 ;
  LAYER M6_m ; RECT -0.5 -0.5 0.5 0.5 ;
END hb_layer_6
VIA hb_layer_7 DEFAULT
  LAYER hb_layer ; RECT -0.25 -0.25 0.25 0.25 ;
  LAYER M7 ; RECT -0.5 -0.25 0.5 0.25 ;
  LAYER M6_m ; RECT -0.25 -0.5 0.25 0.5 ;
END hb_layer_7
VIA hb_layer_8 DEFAULT
  LAYER hb_layer ; RECT -0.25 -0.25 0.25 0.25 ;
  LAYER M7 ; RECT -0.5 -0.25 0.5 0.25 ;
  LAYER M6_m ; RECT -0.5 -0.25 0.5 0.25 ;
END hb_layer_8

VIA VIA56_m Default
  LAYER M5_m ; RECT -0.012 -0.027 0.012 0.027 ;
  LAYER M6_m ; RECT -0.023 -0.016 0.023 0.016 ;
  LAYER V5_m ; RECT -0.012 -0.016 0.012 0.016 ;
END VIA56_m

VIA VIA45_m Default
  LAYER M4_m ; RECT -0.023 -0.012 0.023 0.012 ;
  LAYER M5_m ; RECT -0.012 -0.023 0.012 0.023 ;
  LAYER V4_m ; RECT -0.012 -0.012 0.012 0.012 ;
END VIA45_m

VIA VIA34_m Default
  LAYER M3_m ; RECT -0.009 -0.017 0.009 0.017 ;
  LAYER M4_m ; RECT -0.02 -0.012 0.02 0.012 ;
  LAYER V3_m ; RECT -0.009 -0.012 0.009 0.012 ;
END VIA34_m

VIA VIA23_m Default
  LAYER M2_m ; RECT -0.014 -0.009 0.014 0.009 ;
  LAYER M3_m ; RECT -0.009 -0.014 0.009 0.014 ;
  LAYER V2_m ; RECT -0.009 -0.009 0.009 0.009 ;
END VIA23_m

VIA VIA12_m Default
  LAYER M1_m ; RECT -0.009 -0.011 0.009 0.011 ;
  LAYER M2_m ; RECT -0.014 -0.009 0.014 0.009 ;
  LAYER V1_m ; RECT -0.009 -0.009 0.009 0.009 ;
END VIA12_m

VIA VIA_M1m_M2add DEFAULT
  LAYER M1_m ;   RECT -0.009 -0.011 0.009 0.011 ;
  LAYER M2_add ; RECT -0.014 -0.009 0.014 0.009 ;
  LAYER V1_add ; RECT -0.009 -0.009 0.009 0.009 ;
END VIA_M1m_M2add

VIA VIA_M2add_M3add DEFAULT
  LAYER M2_add ; RECT -0.014 -0.009 0.014 0.009 ;
  LAYER M3_add ; RECT -0.009 -0.014 0.009 0.014 ;
  LAYER V2_add ; RECT -0.009 -0.009 0.009 0.009 ;
END VIA_M2add_M3add

# ======================================================
# 3) VIARULES (after layers & vias)
# ======================================================

VIARULE M7_M6 GENERATE DEFAULT
  LAYER M6 ; ENCLOSURE 0.011 0.0 ;
  LAYER M7 ; ENCLOSURE 0.0 0.011 ;
  LAYER V6 ;
    RECT -0.016 -0.016 0.016 0.016 ;
    SPACING 0.078 BY 0.078 ;
END M7_M6

VIARULE M6_M5 GENERATE DEFAULT
  LAYER M5 ; ENCLOSURE 0.011 0.0 ; WIDTH 0.024 TO 0.024 ;
  LAYER M6 ; ENCLOSURE 0.011 0.0 ; WIDTH 0.032 TO 0.032 ;
  LAYER V5 ;
    RECT -0.012 -0.016 0.012 0.016 ;
    SPACING 0.058 BY 0.308 ; # avoid dual cut on routing
END M6_M5

VIARULE M3_M2widePWR0p936 GENERATE
  LAYER M2 ; ENCLOSURE 0.0 0.0 ;
  LAYER M3 ; ENCLOSURE 0.0 0.0 ; WIDTH 0.234 TO 0.234 ;
  LAYER V2 ;
    RECT -0.117 -0.009 0.117 0.009 ;
    SPACING 0.277 BY 0.036 ;
END M3_M2widePWR0p936

VIARULE M4_M3widePWR0p864 GENERATE
  LAYER M3 ; ENCLOSURE 0.0 0.0 ; WIDTH 0.2335 TO 0.2345 ;
  LAYER M4 ; ENCLOSURE 0.0 0.0 ; WIDTH 0.2155 TO 0.2165 ;
  LAYER V3 ;
    RECT -0.009 -0.108 0.009 0.108 ;
    SPACING 0.036 BY 0.277 ;
END M4_M3widePWR0p864

VIARULE M5_M4widePWR0p864 GENERATE
  LAYER M4 ; ENCLOSURE 0.0 0.0 ;
  LAYER M5 ; ENCLOSURE 0.0 0.0 ; WIDTH 0.216 TO 0.216 ;
  LAYER V4 ;
    RECT -0.108 -0.012 0.108 0.012 ;
    SPACING 0.532 BY 0.096 ;
END M5_M4widePWR0p864

VIARULE M6_M5widePWR1p152 GENERATE
  LAYER M5 ; ENCLOSURE 0.0 0.0 ;
  LAYER M6 ; ENCLOSURE 0.0 0.0 ; WIDTH 0.288 TO 0.288 ;
  LAYER V5 ;
    RECT -0.012 -0.144 0.012 0.144 ;
    SPACING 0.096 BY 0.382 ;
END M6_M5widePWR1p152

VIARULE M7_M6widePWR1p152 GENERATE
  LAYER M6 ; ENCLOSURE 0.0 0.0 ;
  LAYER M7 ; ENCLOSURE 0.0 0.0 ;
  LAYER V6 ;
    RECT -0.144 -0.016 0.144 0.016 ;
    SPACING 0.532 BY 0.096 ;
END M7_M6widePWR1p152

VIARULE M2_M1 GENERATE DEFAULT
  LAYER M1 ; ENCLOSURE 0.0 0.0 ;
  LAYER M2 ; ENCLOSURE 0.002 0.0 ;
  LAYER V1 ;
    RECT -0.009 -0.009 0.009 0.009 ;
    SPACING 0.036 BY 0.036 ;
END M2_M1

VIARULE hb_layerArray-0 GENERATE
  LAYER M7 ;
    ENCLOSURE 0 0 ;
  LAYER M6_m ;
    ENCLOSURE 0 0 ;
  LAYER hb_layer ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1.05 BY 1.05 ;
END hb_layerArray-0

VIARULE M6_m_M5_m GENERATE DEFAULT
  LAYER M5_m ; ENCLOSURE 0.011 0.0 ; WIDTH 0.024 TO 0.024 ;
  LAYER M6_m ; ENCLOSURE 0.011 0.0 ; WIDTH 0.032 TO 0.032 ;
  LAYER V5_m ;
    RECT -0.012 -0.016 0.012 0.016 ;
    SPACING 0.058 BY 0.308 ;
END M6_m_M5_m

VIARULE M3_m_M2_mwidePWR0p936 GENERATE
  LAYER M2_m ; 
    ENCLOSURE 0.0 0.0 ;
  LAYER M3_m ; 
    ENCLOSURE 0.0 0.0 ; WIDTH 0.234 TO 0.234 ;
  LAYER V2_m ;
    RECT -0.117 -0.009 0.117 0.009 ;
    SPACING 0.277 BY 0.036 ;
END M3_m_M2_mwidePWR0p936

VIARULE M4_m_M3_mwidePWR0p864 GENERATE
  LAYER M3_m ; 
    ENCLOSURE 0.0 0.0 ; 
    WIDTH 0.2335 TO 0.2345 ;
  LAYER M4_m ; 
    ENCLOSURE 0.0 0.0 ; 
    WIDTH 0.2155 TO 0.2165 ;
  LAYER V3_m ;
    RECT -0.009 -0.108 0.009 0.108 ;
    SPACING 0.036 BY 0.277 ;
END M4_m_M3_mwidePWR0p864

VIARULE M5_m_M4_mwidePWR0p864 GENERATE
  LAYER M4_m ; ENCLOSURE 0.0 0.0 ;
  LAYER M5_m ; ENCLOSURE 0.0 0.0 ; WIDTH 0.216 TO 0.216 ;
  LAYER V4_m ;
    RECT -0.108 -0.012 0.108 0.012 ;
    SPACING 0.532 BY 0.096 ;
END M5_m_M4_mwidePWR0p864

VIARULE M6_m_M5_mwidePWR1p152 GENERATE
  LAYER M5_m ; ENCLOSURE 0.0 0.0 ;
  LAYER M6_m ; ENCLOSURE 0.0 0.0 ; WIDTH 0.288 TO 0.288 ;
  LAYER V5_m ;
    RECT -0.012 -0.144 0.012 0.144 ;
    SPACING 0.096 BY 0.382 ;
END M6_m_M5_mwidePWR1p152

VIARULE M2_m_M1_m GENERATE DEFAULT
  LAYER M1_m ; ENCLOSURE 0.0 0.0 ;
  LAYER M2_m ; ENCLOSURE 0.002 0.0 ;
  LAYER V1_m ;
    RECT -0.009 -0.009 0.009 0.009 ;
    SPACING 0.036 BY 0.036 ;
END M2_m_M1_m

VIARULE M2add_M1m GENERATE DEFAULT
  LAYER M1_m ; ENCLOSURE 0.0 0.0 ;
  LAYER M2_add ; ENCLOSURE 0.002 0.0 ;
  LAYER V1_add ;
    RECT -0.009 -0.009 0.009 0.009 ;
    SPACING 0.036 BY 0.036 ;
END M2add_M1m

VIARULE M3add_M2add GENERATE DEFAULT
  LAYER M2_add ; ENCLOSURE 0.0 0.0 ;
  LAYER M3_add ; ENCLOSURE 0.0 0.0 ;
  LAYER V2_add ;
    RECT -0.009 -0.009 0.009 0.009 ;
    SPACING 0.036 BY 0.036 ;
END M3add_M2add

END LIBRARY

MACRO HBT_BUF_bottom
  CLASS COVER ;
  ORIGIN 0.0 0.0 ;
  SIZE 0.8 BY 0.8 ;  
  SYMMETRY X Y R90 ;
  SITE CORE ;         

  PIN HB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 0.0 0.0 0.8 0.8 ;
    END
  END HB

END HBT_BUF_bottom

MACRO HBT_BUF_T
  CLASS COVER ;
  ORIGIN 0.0 0.0 ;
  SIZE 0.8 BY 0.8 ;   
  SYMMETRY X Y R90 ;
  SITE CORE ;         

  PIN HB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M6_m ;
        RECT 0.0 0.0 0.8 0.8 ;
    END
  END HB

END HBT_BUF_T
