# BSD 3-Clause License
# 
# Copyright 2020 Lawrence T. Clark, Vinay Vashishtha, or Arizona State
# University
# 
# Redistribution and use in source and binary forms, with or without
# modification, are permitted provided that the following conditions are met:
# 
# 1. Redistributions of source code must retain the above copyright notice,
# this list of conditions and the following disclaimer.
# 
# 2. Redistributions in binary form must reproduce the above copyright
# notice, this list of conditions and the following disclaimer in the
# documentation and/or other materials provided with the distribution.
# 
# 3. Neither the name of the copyright holder nor the names of its
# contributors may be used to endorse or promote products derived from this
# software without specific prior written permission.
# 
# THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
# AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
# IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
# ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
# LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
# CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
# SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
# INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
# CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
# ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
# POSSIBILITY OF SUCH DAMAGE.

VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
CLEARANCEMEASURE EUCLIDEAN ;
USEMINSPACING OBS OFF ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.001 ;

# ========================
# Property Definitions
# ========================
PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_PITCH STRING ;
  LAYER LEF58_GAP STRING ;
  LAYER LEF58_EOLKEEPOUT STRING ;
  LAYER LEF58_SPACING STRING ;
  LAYER LEF58_CORNERSPACING STRING ;
  LAYER LEF58_WIDTHTABLE STRING ;
  LAYER LEF58_CUTCLASS STRING ;
  LAYER LEF58_SPACINGTABLE STRING ;
  LAYER LEF58_ENCLOSURE STRING ;
  LAYER LEF58_RIGHTWAYONGRIDONLY STRING ;
  LAYER LEF58_RECTONLY STRING ;
END PROPERTYDEFINITIONS

LAYER nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END pwell

LAYER poly
  TYPE MASTERSLICE ;
END poly

LAYER active
  TYPE MASTERSLICE ;
END active

LAYER M1
  TYPE ROUTING ;
  SPACING 0.065 ;
  WIDTH 0.07 ;
  PITCH 0.14 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.38 ;
  THICKNESS 0.13 ;
  HEIGHT 0.37 ;
  CAPACITANCE CPERSQDIST 7.7161e-05 ;
  EDGECAPACITANCE 2.7365e-05 ;
END M1

LAYER via1
  TYPE CUT ;
  SPACING 0.08 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via1

LAYER M2
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.3000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.0700     0.0700     0.0700     0.0700     0.0700     0.0700     
      WIDTH 0.0900       0.0700     0.0900     0.0900     0.0900     0.0900     0.0900     
      WIDTH 0.2700       0.0700     0.0900     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.0700     0.0900     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.0700     0.0900     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.0700     0.0900     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.07 ;
  PITCH 0.19 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  HEIGHT 0.62 ;
  CAPACITANCE CPERSQDIST 4.0896e-05 ;
  EDGECAPACITANCE 2.5157e-05 ;
END M2

LAYER via2
  TYPE CUT ;
  SPACING 0.09 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via2

LAYER M3
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.3000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.0700     0.0700     0.0700     0.0700     0.0700     0.0700     
      WIDTH 0.0900       0.0700     0.0900     0.0900     0.0900     0.0900     0.0900     
      WIDTH 0.2700       0.0700     0.0900     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.0700     0.0900     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.0700     0.0900     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.0700     0.0900     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.07 ;
  PITCH 0.14 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  HEIGHT 0.88 ;
  CAPACITANCE CPERSQDIST 2.7745e-05 ;
  EDGECAPACITANCE 2.5157e-05 ;
END M3

LAYER via3
  TYPE CUT ;
  SPACING 0.09 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via3

LAYER M4
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400     
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 1.14 ;
  CAPACITANCE CPERSQDIST 2.0743e-05 ;
  EDGECAPACITANCE 3.0908e-05 ;
END M4

LAYER via4
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via4

LAYER M5
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400     
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 1.71 ;
  CAPACITANCE CPERSQDIST 1.3527e-05 ;
  EDGECAPACITANCE 2.3863e-06 ;
END M5

LAYER via5
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via5

LAYER M6
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400     
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 2.28 ;
  CAPACITANCE CPERSQDIST 1.0036e-05 ;
  EDGECAPACITANCE 2.3863e-05 ;
END M6

LAYER via6
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via6

LAYER M7
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.4000     0.4000     0.4000     0.4000     
      WIDTH 0.5000       0.4000     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.4000     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.4000     0.5000     0.9000     1.5000      ;
  WIDTH 0.4 ;
  PITCH 0.8 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.075 ;
  THICKNESS 0.8 ;
  HEIGHT 2.85 ;
  CAPACITANCE CPERSQDIST 7.9771e-06 ;
  EDGECAPACITANCE 3.2577e-05 ;
END M7

LAYER via7
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  RESISTANCE 1 ;
END via7

LAYER M8
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.4000     0.4000     0.4000     0.4000     
      WIDTH 0.5000       0.4000     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.4000     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.4000     0.5000     0.9000     1.5000      ;
  WIDTH 0.4 ;
  PITCH 0.8 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.075 ;
  THICKNESS 0.8 ;
  HEIGHT 4.47 ;
  CAPACITANCE CPERSQDIST 5.0391e-06 ;
  EDGECAPACITANCE 2.3932e-05 ;
END M8

LAYER via8
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  RESISTANCE 1 ;
END via8

LAYER M9
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     2.7000     4.0000     
      WIDTH 0.0000       0.8000     0.8000     0.8000     
      WIDTH 0.9000       0.8000     0.9000     0.9000     
      WIDTH 1.5000       0.8000     0.9000     1.5000      ;
  WIDTH 0.8 ;
  PITCH 1.6 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.03 ;
  THICKNESS 2 ;
  HEIGHT 6.09 ;
  CAPACITANCE CPERSQDIST 3.6827e-06 ;
  EDGECAPACITANCE 3.0803e-05 ;
END M9

LAYER via9
  TYPE CUT ;
  SPACING 0.88 ;
  WIDTH 0.8 ;
  RESISTANCE 0.5 ;
END via9

LAYER M10
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     2.7000     4.0000     
      WIDTH 0.0000       0.8000     0.8000     0.8000     
      WIDTH 0.9000       0.8000     0.9000     0.9000     
      WIDTH 1.5000       0.8000     0.9000     1.5000      ;
  WIDTH 0.8 ;
  PITCH 1.6 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.03 ;
  THICKNESS 2 ;
  HEIGHT 10.09 ;
  CAPACITANCE CPERSQDIST 2.2124e-06 ;
  EDGECAPACITANCE 2.3667e-05 ;
END M10

LAYER hb_layer
  TYPE CUT ;
  SPACING 0.8 ;
  WIDTH 0.8 ;
  RESISTANCE 0.02 ;
END hb_layer

LAYER M8_m
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.08 0.08 ;
  WIDTH 0.04 ;
  AREA 0.00752 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0 0.39975 1.19975 1.79975
    WIDTH 0.0 0.04 0.04 0.04 0.04
    WIDTH 0.05975 0.04 0.04 0.04 0.04
    WIDTH 0.07975 0.04 0.04 0.04 0.04
    WIDTH 0.11975 0.04 0.04 0.04 0.04
    WIDTH 0.49975 0.04 0.04 0.04 0.5
    WIDTH 0.99975 0.04 0.04 0.04 1.0 ;
  MINIMUMCUT 2 WIDTH 1.805 WITHIN 1.705 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 1.805 WITHIN 1.705 FROMABOVE ;
  MAXWIDTH 2.0 ;
  MINSTEP 0.04 STEP ;
# --- RC added from ict/setRC for M8_m ---
  THICKNESS 0.08 ;
  HEIGHT 12.41 ;
  RESISTANCE RPERSQ 0.474476 ;
  CAPACITANCE CPERSQDIST 0.001321 ;
  EDGECAPACITANCE 6.165110e-05 ;
END M8_m

LAYER V7_m
  TYPE CUT ;
  SPACING 0.046 ;
  WIDTH 0.032 ;
# --- RC added from ict/setRC for V7_m ---
  RESISTANCE 8.2 ;
END V7_m

LAYER M7_m
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.064 ;
  WIDTH 0.032 ;
  SPACING 0.032 ;
  AREA 0.0021875 ;
  PROPERTY LEF58_SPACING " SPACING 0.03 ENDOFLINE 0.0375 WITHIN 0.04 ENDTOEND 0.04 ; " ;
  PROPERTY LEF58_WIDTHTABLE " WIDTHTABLE 0.032 0.16 0.288 0.416 0.544 ; " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER CORNERONLY 0.075
   WIDTH 0.0 SPACING 0.04 ;
   " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.05 EXTENSION 0.048 0.03225 0.048
      CORNERONLY ;
   " ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0
    WIDTH 0.0 0.032
    WIDTH 0.033 0.072 ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M7_m ---
  THICKNESS 0.064 ;
  HEIGHT 12.538 ;
  RESISTANCE RPERSQ 0.400995 ;
  CAPACITANCE CPERSQDIST 0.001378 ;
  EDGECAPACITANCE 5.146050e-05 ;
END M7_m

LAYER V6_m
  TYPE CUT ;
  PROPERTY LEF58_CUTCLASS "
   CUTCLASS Vx WIDTH 0.032 LENGTH 0.032 ;
   CUTCLASS Vx_0p640 WIDTH 0.032 LENGTH 0.16 CUTS 4 ;
   CUTCLASS Vx_1p152 WIDTH 0.032 LENGTH 0.288 CUTS 8 ;
   CUTCLASS Vx_1p664 WIDTH 0.032 LENGTH 0.416 CUTS 12 ;
   CUTCLASS Vx_2p176 WIDTH 0.032 LENGTH 0.544 CUTS 16 ;
   " ;
  PROPERTY LEF58_SPACINGTABLE "
      SPACINGTABLE
       DEFAULT 0.034
       CUTCLASS Vx Vx_0p640 Vx_1p152 Vx_1p664 Vx_2p176
              Vx       -  -        -        -        - -  -        -        -        -
              Vx_0p640 -  -        -        -        - -  -        -        -        -
	      Vx_1p152 -  -        -        -        - -  -        -        -        -
	      Vx_1p664 -  -        -        -        - -  -        -        -        -
	      Vx_2p176 -  -        -        -        - -  -        -        -        -
      ;
   " ;
  PROPERTY LEF58_ENCLOSURE "
   ENCLOSURE CUTCLASS Vx 0.011 0.0 ;
   ENCLOSURE CUTCLASS Vx EOL 0.0 0.011 0.011 ;
   ENCLOSURE CUTCLASS Vx_0p640 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p152 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p664 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_2p176 END 0.0 SIDE 0.0 ;
   " ;
# --- RC added from ict/setRC for V6_m ---
  RESISTANCE 8.2 ;
END V6_m

LAYER M6_m
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.064 ;
  WIDTH 0.032 ;
  SPACING 0.032 ;
  AREA 0.0021875 ;
  PROPERTY LEF58_SPACING " SPACING 0.032 ENDOFLINE 0.0375 WITHIN 0.04 ENDTOEND 0.04 ; " ;
  PROPERTY LEF58_WIDTHTABLE " WIDTHTABLE 0.032 0.16 0.288 0.416 0.544 ; " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER CORNERONLY 0.048
   WIDTH 0.0 SPACING 0.04 ;
   " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.05 EXTENSION 0.048 0.03225 0.048 CORNERONLY ;
   " ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0
    WIDTH 0.0 0.032
    WIDTH 0.033 0.072 ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M6_m ---
  THICKNESS 0.064 ;
  HEIGHT 12.666 ;
  RESISTANCE RPERSQ 0.379581 ;
  CAPACITANCE CPERSQDIST 0.001651 ;
  EDGECAPACITANCE 6.165110e-05 ;
END M6_m

LAYER V5_m
  TYPE CUT ;
  PROPERTY LEF58_CUTCLASS "
   CUTCLASS Vx WIDTH 0.024 LENGTH 0.032 ;
   CUTCLASS Vx_0p480 WIDTH 0.024 LENGTH 0.16 CUTS 4 ;
   CUTCLASS Vx_0p864 WIDTH 0.024 LENGTH 0.288 CUTS 8 ;
   CUTCLASS Vx_1p248 WIDTH 0.024 LENGTH 0.416 CUTS 12 ;
   CUTCLASS Vx_1p632 WIDTH 0.024 LENGTH 0.544 CUTS 16 ;
   " ;
  PROPERTY LEF58_SPACINGTABLE "
      SPACINGTABLE
       DEFAULT 0.034
       CUTCLASS Vx Vx_0p480 Vx_0p864 Vx_1p248 Vx_1p632
              Vx       -  -        -        -        - -  -        -        -        -
              Vx_0p480 -  -        -        -        - -  -        -        -        -
	      Vx_0p864 -  -        -        -        - -  -        -        -        -
	      Vx_1p248 -  -        -        -        - -  -        -        -        -
	      Vx_1p632 -  -        -        -        - -  -        -        -        -
      ;
   " ;
  PROPERTY LEF58_ENCLOSURE "
   ENCLOSURE CUTCLASS Vx EOL 0.02425 0.011 0.011 ;
   ENCLOSURE CUTCLASS Vx_0p480 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_0p864 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p248 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p632 END 0.0 SIDE 0.0 ;
   " ;
# --- RC added from ict/setRC for V5_m ---
  RESISTANCE 11.8 ;
END V5_m

LAYER M5_m
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.048 ;
  WIDTH 0.024 ;
  SPACING 0.024 ;
  OFFSET 0.0 ;
  AREA 0.002 ;
  PROPERTY LEF58_SPACING " SPACING 0.024 ENDOFLINE 0.025 WITHIN 0.04 ENDTOEND 0.04 ; " ;
  MINIMUMDENSITY 15.0 ;
  MAXIMUMDENSITY 90.0 ;
  DENSITYCHECKWINDOW 20.0 20.0 ;
  DENSITYCHECKSTEP 10.0 ;
  PROPERTY LEF58_WIDTHTABLE
   " WIDTHTABLE 0.024 0.12 0.216 0.312 0.408 0.504 0.6 0.696 0.792 0.888 0.984 ; " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER CORNERONLY 0.048
   WIDTH 0.0 SPACING 0.04 ;
   " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.025 EXTENSION 0.048 0.02425 0.048
      CORNERONLY ;
   " ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0
    WIDTH 0.0 0.024
    WIDTH 0.025 0.072 ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M5_m ---
  THICKNESS 0.048 ;
  HEIGHT 12.762 ;
  RESISTANCE RPERSQ 0.463212 ;
  CAPACITANCE CPERSQDIST 0.002145 ;
  EDGECAPACITANCE 6.005755e-05 ;
END M5_m

LAYER V4_m
  TYPE CUT ;
  PROPERTY LEF58_CUTCLASS "
   CUTCLASS Vx WIDTH 0.024 LENGTH 0.024 ;
   CUTCLASS Vx_0p480 WIDTH 0.024 LENGTH 0.12 CUTS 4 ;
   CUTCLASS Vx_0p864 WIDTH 0.024 LENGTH 0.216 CUTS 8 ;
   CUTCLASS Vx_1p248 WIDTH 0.024 LENGTH 0.312 CUTS 12 ;
   CUTCLASS Vx_1p632 WIDTH 0.024 LENGTH 0.408 CUTS 16 ;
   " ;
  PROPERTY LEF58_SPACINGTABLE "
      SPACINGTABLE
       DEFAULT 0.034
       CUTCLASS Vx Vx_0p480 Vx_0p864 Vx_1p248 Vx_1p632
              Vx       -  -        -        -        - -  -        -        -        -
              Vx_0p480 -  -        -        -        - -  -        -        -        -
	      Vx_0p864 -  -        -        -        - -  -        -        -        -
	      Vx_1p248 -  -        -        -        - -  -        -        -        -
	      Vx_1p632 -  -        -        -        - -  -        -        -        -
      ;
   " ;
  PROPERTY LEF58_ENCLOSURE "
   ENCLOSURE CUTCLASS Vx 0.011 0.0 ;
   ENCLOSURE CUTCLASS Vx EOL 0.0 0.011 0.011 ;
   ENCLOSURE CUTCLASS Vx_0p480 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_0p864 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p248 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS Vx_1p632 END 0.0 SIDE 0.0 ;
   " ;
# --- RC added from ict/setRC for V4_m ---
  RESISTANCE 11.8 ;
END V4_m

LAYER M4_m
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.048 ;
  WIDTH 0.024 ;
  SPACING 0.024 ;
  OFFSET 0.003 ;
  AREA 0.002 ;
  PROPERTY LEF58_SPACING " SPACING 0.024 ENDOFLINE 0.025 WITHIN 0.04 ENDTOEND 0.04 ; " ;
  PROPERTY LEF58_WIDTHTABLE " WIDTHTABLE 0.024 0.12 0.216 0.312 0.408 ; " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER CORNERONLY 0.048
   WIDTH 0.0 SPACING 0.04 ;
   " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.025 EXTENSION 0.048 0.02425 0.048 CORNERONLY ;
   " ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0
    WIDTH 0.0 0.024
    WIDTH 0.025 0.072 ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M4_m ---
  THICKNESS 0.048 ;
  HEIGHT 12.858 ;
  RESISTANCE RPERSQ 0.487399 ;
  CAPACITANCE CPERSQDIST 0.002368 ;
  EDGECAPACITANCE 6.630190e-05 ;
END M4_m

LAYER V3_m
  TYPE CUT ;
  PROPERTY LEF58_CUTCLASS "
   CUTCLASS V3 WIDTH 0.018 LENGTH 0.024 CUTS 1 ;
   CUTCLASS V3_0p480 WIDTH 0.018 LENGTH 0.12 CUTS 4 ;
   CUTCLASS V3_0p864 WIDTH 0.018 LENGTH 0.216 CUTS 8 ;
   " ;
  PROPERTY LEF58_SPACINGTABLE "
      SPACINGTABLE
       DEFAULT 0.034
       CUTCLASS V3 V3_0p480 V3_0p864
              V3       -  -        -        -  - -
              V3_0p480 -  -        -        -  - -
              V3_0p864 -  -        -        -  - -
      ;
   " ;
  PROPERTY LEF58_ENCLOSURE "
   ENCLOSURE CUTCLASS V3 BELOW EOL 0.0 0.005 0.0 ;
   ENCLOSURE CUTCLASS V3 ABOVE EOL 0.02425 0.011 0.0 ;
   ENCLOSURE CUTCLASS V3_0p480 END 0.0 SIDE 0.0 ;
   ENCLOSURE CUTCLASS V3_0p864 END 0.0 SIDE 0.0 ;
   " ;
# --- RC added from ict/setRC for V3_m ---
  RESISTANCE 17.2 ;
END V3_m

LAYER M3_m
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.036 ;
  OFFSET 0.0 ;
  WIDTH 0.018 ;
  SPACING 0.018 ;
  AREA 0.000666 ;
  MINSIZE 0.037 0.018 ;
  PROPERTY LEF58_SPACING
   " SPACING 0.018 ENDOFLINE 0.025 WITHIN 0.0125 ENDTOEND 0.031
     PARALLELEDGE 0.025 WITHIN 0.02 ; " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.025 EXTENSION 0.0 0.0125 0.031 CORNERONLY ;
   " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER WIDTH 0.0 SPACING 0.02
     ;
   " ;
  PROPERTY LEF58_WIDTHTABLE
   " WIDTHTABLE 0.018 0.09 0.162 0.234 0.306 0.378 ; " ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M3_m ---
  THICKNESS 0.036 ;
  HEIGHT 12.93 ;
  RESISTANCE RPERSQ 0.653852 ;
  CAPACITANCE CPERSQDIST 0.002566 ;
  EDGECAPACITANCE 5.388425e-05 ;
END M3_m

LAYER V2_m
  TYPE CUT ;
  SPACING 0.018 ;
  WIDTH 0.018 ;
# --- RC added from ict/setRC for V2_m ---
  RESISTANCE 17.2 ;
END V2_m

LAYER M2_m
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.018 ;
  SPACING 0.018 ;
  OFFSET -0.27 ;
  AREA 0.000666 ;
  MINSIZE 0.037 0.018 ;
  PITCH 0.045 0.036 ;
  PROPERTY LEF58_PITCH "
   PITCH 0.036 FIRSTLASTPITCH 0.045
     ;
   " ;
  PROPERTY LEF58_SPACING
   " SPACING 0.018 ENDOFLINE 0.025 WITHIN 0.02 ENDTOEND 0.031
     PARALLELEDGE 0.025 WITHIN 0.02 ; " ;
  PROPERTY LEF58_EOLKEEPOUT "
   EOLKEEPOUT 0.025 EXTENSION 0.0 0.0125 0.031 CORNERONLY ;
   " ;
  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER WIDTH 0.0 SPACING 0.02 ;
   " ;
  PROPERTY LEF58_WIDTHTABLE "
   WIDTHTABLE 0.018 0.09 0.162 0.234 0.306 0.378 ;
   " ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY " RIGHTWAYONGRIDONLY ; " ;
  PROPERTY LEF58_RECTONLY " RECTONLY ; " ;
# --- RC added from ict/setRC for M2_m ---
  THICKNESS 0.036 ;
  HEIGHT 13.002 ;
  RESISTANCE RPERSQ 0.83216 ;
  CAPACITANCE CPERSQDIST 0.003076 ;
  EDGECAPACITANCE 6.458970e-05 ;
END M2_m

LAYER V1_m
  TYPE CUT ;
  SPACING 0.018 ;
  WIDTH 0.018 ;
# --- RC added from ict/setRC for V1_m ---
  RESISTANCE 17.2 ;
END V1_m

LAYER M1_m
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.036 ;
  WIDTH 0.018 ;
  SPACING 0.018 ;
  AREA 0.000666 ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.01825 EXTENSION 0.0 0.0 0.031 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERONLY 0.01 WIDTH 0.018 SPACING 0.018 ;" ;
  OFFSET 0.0 ;
# --- RC added from ict/setRC for M1_m ---
  THICKNESS 0.036 ;
  HEIGHT 13.074 ;
  RESISTANCE RPERSQ 1.267515 ;
  CAPACITANCE CPERSQDIST 1.000000e-08 ;
  EDGECAPACITANCE 1.000000e-08 ;
END M1_m

# LAYER V0_m
#   TYPE CUT ;
#   SPACING 0.018 ;
#   WIDTH 0.018 ;
# END V0_m

LAYER RVTN_m
  TYPE IMPLANT ;
END RVTN_m

LAYER RVTP_m
  TYPE IMPLANT ;
END RVTP_m

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

# ======================================================
# 2) VIA MACROS (after all layers)
# ======================================================

VIA via1_4 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via1_4

VIA via1_0 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1_0

VIA via1_1 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via1_1

VIA via1_2 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via1_2

VIA via1_3 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1_3

VIA via1_5 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via1_5

VIA via1_6 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1_6

VIA via1_7 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via1_7

VIA via1_8 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via1_8

VIA via2_8 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via2_8

VIA via2_4 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via2_4

VIA via2_5 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via2_5

VIA via2_7 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via2_7

VIA via2_6 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2_6

VIA via2_0 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2_0

VIA via2_1 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via2_1

VIA via2_2 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via2_2

VIA via2_3 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2_3

VIA via3_2 DEFAULT
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3_2

VIA via3_0 DEFAULT
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3_0

VIA via3_1 DEFAULT
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER M3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3_1

VIA via4_0 DEFAULT
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via4_0

VIA via5_0 DEFAULT
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via5_0

VIA via6_0 DEFAULT
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER M7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END via6_0

VIA via7_0 DEFAULT
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER M7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER M8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END via7_0

VIA via8_0 DEFAULT
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER M8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER M9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END via8_0

VIA via9_0 DEFAULT
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER M9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER M10 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END via9_0

VIA hb_layer_0 DEFAULT
  LAYER hb_layer ; RECT -0.4 -0.4 0.4 0.4 ;
  LAYER M10 ; RECT -0.4 -0.4 0.4 0.4 ;
  LAYER M8_m ; RECT -0.4 -0.4 0.4 0.4 ;
END hb_layer_0

VIA hb_layer_1 DEFAULT
  LAYER hb_layer ; RECT -0.4 -0.4 0.4 0.4 ;
  LAYER M10 ; RECT -0.8 -0.8 0.8 0.8 ;
  LAYER M8_m ; RECT -0.4 -0.8 0.4 0.8 ;
END hb_layer_1

VIA hb_layer_2 DEFAULT
  LAYER hb_layer ; RECT -0.4 -0.4 0.4 0.4 ;
  LAYER M10 ; RECT -0.8 -0.8 0.8 0.8 ;
  LAYER M8_m ; RECT -0.8 -0.4 0.8 0.4 ;
END hb_layer_2

VIA hb_layer_3 DEFAULT
  LAYER hb_layer ; RECT -0.4 -0.4 0.4 0.4 ;
  LAYER M10 ; RECT -0.4 -0.8 0.4 0.8 ;
  LAYER M8_m ; RECT -0.8 -0.8 0.8 0.8 ;
END hb_layer_3

VIA hb_layer_4 DEFAULT
  LAYER hb_layer ; RECT -0.4 -0.4 0.4 0.4 ;
  LAYER M10 ; RECT -0.4 -0.8 0.4 0.8 ;
  LAYER M8_m ; RECT -0.4 -0.8 0.4 0.8 ;
END hb_layer_4

VIA hb_layer_5 DEFAULT
  LAYER hb_layer ; RECT -0.4 -0.4 0.4 0.4 ;
  LAYER M10 ; RECT -0.4 -0.8 0.4 0.8 ;
  LAYER M8_m ; RECT -0.8 -0.4 0.8 0.4 ;
END hb_layer_5

VIA hb_layer_6 DEFAULT
  LAYER hb_layer ; RECT -0.4 -0.4 0.4 0.4 ;
  LAYER M10 ; RECT -0.8 -0.4 0.8 0.4 ;
  LAYER M8_m ; RECT -0.8 -0.8 0.8 0.8 ;
END hb_layer_6

VIA hb_layer_7 DEFAULT
  LAYER hb_layer ; RECT -0.4 -0.4 0.4 0.4 ;
  LAYER M10 ; RECT -0.8 -0.4 0.8 0.4 ;
  LAYER M8_m ; RECT -0.4 -0.8 0.4 0.8 ;
END hb_layer_7

VIA hb_layer_8 DEFAULT
  LAYER hb_layer ; RECT -0.4 -0.4 0.4 0.4 ;
  LAYER M10 ; RECT -0.8 -0.4 0.8 0.4 ;
  LAYER M8_m ; RECT -0.8 -0.4 0.8 0.4 ;
END hb_layer_8

VIA VIA12_m Default
  LAYER M1_m ; RECT -0.009 -0.011 0.009 0.011 ;
  LAYER M2_m ; RECT -0.014 -0.009 0.014 0.009 ;
  LAYER V1_m ; RECT -0.009 -0.009 0.009 0.009 ;
END VIA12_m

VIA VIA23_m Default
  LAYER M2_m ; RECT -0.014 -0.009 0.014 0.009 ;
  LAYER M3_m ; RECT -0.009 -0.014 0.009 0.014 ;
  LAYER V2_m ; RECT -0.009 -0.009 0.009 0.009 ;
END VIA23_m

VIA VIA34_m Default
  LAYER M3_m ; RECT -0.009 -0.017 0.009 0.017 ;
  LAYER M4_m ; RECT -0.02 -0.012 0.02 0.012 ;
  LAYER V3_m ; RECT -0.009 -0.012 0.009 0.012 ;
END VIA34_m

VIA VIA45_m Default
  LAYER M4_m ; RECT -0.023 -0.012 0.023 0.012 ;
  LAYER M5_m ; RECT -0.012 -0.023 0.012 0.023 ;
  LAYER V4_m ; RECT -0.012 -0.012 0.012 0.012 ;
END VIA45_m

VIA VIA56_m Default
  LAYER M5_m ; RECT -0.012 -0.027 0.012 0.027 ;
  LAYER M6_m ; RECT -0.023 -0.016 0.023 0.016 ;
  LAYER V5_m ; RECT -0.012 -0.016 0.012 0.016 ;
END VIA56_m

VIA VIA67_m Default
  LAYER M6_m ; RECT -0.027 -0.016 0.027 0.016 ;
  LAYER M7_m ; RECT -0.016 -0.027 0.016 0.027 ;
  LAYER V6_m ; RECT -0.016 -0.016 0.016 0.016 ;
END VIA67_m

VIA VIA78_m Default
  LAYER M7_m ; RECT -0.016 -0.027 0.016 0.027 ;
  LAYER M8_m ; RECT -0.027 -0.020 0.027 0.020 ;
  LAYER V7_m ; RECT -0.016 -0.016 0.016 0.016 ;
END VIA78_m

# ======================================================
# 3) VIARULES (after layers & vias)
# ======================================================

VIARULE M8_m_M7_m GENERATE DEFAULT
  LAYER M7_m ; ENCLOSURE 0.0 0.0 ;
  LAYER M8_m ; ENCLOSURE 0.011 0.0 ;
  LAYER V7_m ;
    RECT -0.016 -0.016 0.016 0.016 ;
    SPACING 0.078 BY 0.078 ;
END M8_m_M7_m

VIARULE M7_m_M6_m GENERATE DEFAULT
  LAYER M6_m ; ENCLOSURE 0.011 0.0 ;
  LAYER M7_m ; ENCLOSURE 0.0 0.011 ;
  LAYER V6_m ;
    RECT -0.016 -0.016 0.016 0.016 ;
    SPACING 0.078 BY 0.078 ;
END M7_m_M6_m

VIARULE M6_m_M5_m GENERATE DEFAULT
  LAYER M5_m ; ENCLOSURE 0.011 0.0 ; WIDTH 0.024 TO 0.024 ;
  LAYER M6_m ; ENCLOSURE 0.011 0.0 ; WIDTH 0.032 TO 0.032 ;
  LAYER V5_m ;
    RECT -0.012 -0.016 0.012 0.016 ;
    SPACING 0.058 BY 0.308 ;
END M6_m_M5_m


VIARULE M3_m_M2_mwidePWR0p936 GENERATE
  LAYER M2_m ; ENCLOSURE 0.0 0.0 ;
  LAYER M3_m ; ENCLOSURE 0.0 0.0 ; WIDTH 0.234 TO 0.234 ;
  LAYER V2_m ;
    RECT -0.117 -0.009 0.117 0.009 ;
    SPACING 0.277 BY 0.036 ;
END M3_m_M2_mwidePWR0p936

VIARULE M4_m_M3_mwidePWR0p864 GENERATE
  LAYER M3_m ; ENCLOSURE 0.0 0.0 ; WIDTH 0.2335 TO 0.2345 ;
  LAYER M4_m ; ENCLOSURE 0.0 0.0 ; WIDTH 0.2155 TO 0.2165 ;
  LAYER V3_m ;
    RECT -0.009 -0.108 0.009 0.108 ;
    SPACING 0.036 BY 0.277 ;
END M4_m_M3_mwidePWR0p864

VIARULE M5_m_M4_mwidePWR0p864 GENERATE
  LAYER M4_m ; ENCLOSURE 0.0 0.0 ;
  LAYER M5_m ; ENCLOSURE 0.0 0.0 ; WIDTH 0.216 TO 0.216 ;
  LAYER V4_m ;
    RECT -0.108 -0.012 0.108 0.012 ;
    SPACING 0.532 BY 0.096 ;
END M5_m_M4_mwidePWR0p864

VIARULE M6_m_M5_mwidePWR1p152 GENERATE
  LAYER M5_m ; ENCLOSURE 0.0 0.0 ;
  LAYER M6_m ; ENCLOSURE 0.0 0.0 ; WIDTH 0.288 TO 0.288 ;
  LAYER V5_m ;
    RECT -0.012 -0.144 0.012 0.144 ;
    SPACING 0.096 BY 0.382 ;
END M6_m_M5_mwidePWR1p152

VIARULE M7_m_M6_mwidePWR1p152 GENERATE
  LAYER M6_m ; ENCLOSURE 0.0 0.0 ;
  LAYER M7_m ; ENCLOSURE 0.0 0.0 ;
  LAYER V6_m ;
    RECT -0.144 -0.016 0.144 0.016 ;
    SPACING 0.532 BY 0.096 ;
END M7_m_M6_mwidePWR1p152

VIARULE M2_m_M1_m GENERATE DEFAULT
  LAYER M1_m ; ENCLOSURE 0.0 0.0 ;
  LAYER M2_m ; ENCLOSURE 0.002 0.0 ;
  LAYER V1_m ;
    RECT -0.009 -0.009 0.009 0.009 ;
    SPACING 0.036 BY 0.036 ;
END M2_m_M1_m

VIARULE hb_layerArray-0 GENERATE
  LAYER M8_m ; ENCLOSURE 0 0 ;
  LAYER M10  ; ENCLOSURE 0 0 ;
  LAYER hb_layer ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 0.4 BY 0.4 ;
END hb_layerArray-0

VIARULE Via1Array-0 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER M2 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-0

VIARULE Via1Array-1 GENERATE
  LAYER M1 ;
    ENCLOSURE 0 0.035 ;
  LAYER M2 ;
    ENCLOSURE 0 0.035 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-1

VIARULE Via1Array-2 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.035 0 ;
  LAYER M2 ;
    ENCLOSURE 0.035 0 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-2

VIARULE Via1Array-3 GENERATE
  LAYER M1 ;
    ENCLOSURE 0 0.035 ;
  LAYER M2 ;
    ENCLOSURE 0.035 0 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-3

VIARULE Via1Array-4 GENERATE
  LAYER M1 ;
    ENCLOSURE 0.035 0 ;
  LAYER M2 ;
    ENCLOSURE 0 0.035 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-4

VIARULE Via2Array-0 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER M3 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-0

VIARULE Via2Array-1 GENERATE
  LAYER M2 ;
    ENCLOSURE 0 0.035 ;
  LAYER M3 ;
    ENCLOSURE 0 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-1

VIARULE Via2Array-2 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.035 0 ;
  LAYER M3 ;
    ENCLOSURE 0.035 0 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-2

VIARULE Via2Array-3 GENERATE
  LAYER M2 ;
    ENCLOSURE 0 0.035 ;
  LAYER M3 ;
    ENCLOSURE 0.035 0 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-3

VIARULE Via2Array-4 GENERATE
  LAYER M2 ;
    ENCLOSURE 0.035 0 ;
  LAYER M3 ;
    ENCLOSURE 0 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-4

VIARULE Via3Array-0 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER M4 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via3Array-0

VIARULE Via3Array-1 GENERATE
  LAYER M3 ;
    ENCLOSURE 0 0.035 ;
  LAYER M4 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via3Array-1

VIARULE Via3Array-2 GENERATE
  LAYER M3 ;
    ENCLOSURE 0.035 0 ;
  LAYER M4 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via3Array-2

VIARULE Via4Array-0 GENERATE
  LAYER M4 ;
    ENCLOSURE 0 0 ;
  LAYER M5 ;
    ENCLOSURE 0 0 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via4Array-0

VIARULE Via5Array-0 GENERATE
  LAYER M5 ;
    ENCLOSURE 0 0 ;
  LAYER M6 ;
    ENCLOSURE 0 0 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via5Array-0

VIARULE Via6Array-0 GENERATE
  LAYER M6 ;
    ENCLOSURE 0 0 ;
  LAYER M7 ;
    ENCLOSURE 0.13 0.13 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via6Array-0

VIARULE Via7Array-0 GENERATE
  LAYER M7 ;
    ENCLOSURE 0 0 ;
  LAYER M8 ;
    ENCLOSURE 0 0 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via7Array-0

VIARULE Via8Array-0 GENERATE
  LAYER M8 ;
    ENCLOSURE 0 0 ;
  LAYER M9 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via8Array-0

VIARULE Via9Array-0 GENERATE
  LAYER M10 ;
    ENCLOSURE 0 0 ;
  LAYER M9 ;
    ENCLOSURE 0 0 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.68 BY 1.68 ;
END Via9Array-0

SPACING
  SAMENET M1 M1 0.065 ;
  SAMENET M2 M2 0.07 ;
  SAMENET M3 M3 0.07 ;
  SAMENET M4 M4 0.14 ;
  SAMENET M5 M5 0.14 ;
  SAMENET M6 M6 0.14 ;
  SAMENET M7 M7 0.4 ;
  SAMENET M8 M8 0.4 ;
  SAMENET M9 M9 0.8 ;
  SAMENET M10 M10 0.8 ;
  SAMENET via1 via1 0.08 ;
  SAMENET via2 via2 0.09 ;
  SAMENET via3 via3 0.09 ;
  SAMENET via4 via4 0.16 ;
  SAMENET via5 via5 0.16 ;
  SAMENET via6 via6 0.16 ;
  SAMENET via7 via7 0.44 ;
  SAMENET via8 via8 0.44 ;
  SAMENET via9 via9 0.88 ;
  SAMENET via1 via2 0.0 STACK ;
  SAMENET via2 via3 0.0 STACK ;
  SAMENET via3 via4 0.0 STACK ;
  SAMENET via4 via5 0.0 STACK ;
  SAMENET via5 via6 0.0 STACK ;
  SAMENET via6 via7 0.0 STACK ;
  SAMENET via7 via8 0.0 STACK ;
  SAMENET via8 via9 0.0 STACK ;
END SPACING

END LIBRARY